`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01.09.2025 10:56:59
// Design Name: 
// Module Name: qns_no_2_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module qns_no_2_tb();
   reg clk, reset, x;
    wire y;

    qns_no_2 uut (
        .clk(clk),
        .reset(reset),
        .x(x),
        .y(y)
    );

    always #5 clk = ~clk;

    reg [15:0] test_vec;
    integer i;

    initial begin
        clk = 0; reset = 1; x = 0;
        #12 reset = 0;
        test_vec = 16'b0101101111010100;
        for (i = 15; i >= 0; i = i - 1) begin
            x = test_vec[i];
            #10;
        end
        #20 $finish;
    end

endmodule

